
module sdc_dsp_core
	(input logic clk,
	 input logic rst);
	 


endmodule
